package agnt_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "agnt1_seq_item.sv"
`include "agnt1_driver.sv"
`include "agnt1_mon.sv"
`include "agnt1_seqr.sv"
`include "agnt1_agent.sv"
`include "agnt2_seq_item.sv"
`include "agnt2_driver.sv"
`include "agnt2_mon.sv"
`include "agnt2_seqr.sv"
`include "agnt2_agent.sv"
endpackage
