interface agnt_name_intf;

    // Declare Struct handles


endinterface
