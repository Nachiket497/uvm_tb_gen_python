package agnt1_pkg;
`include agnt1_seq_item.sv
`include agnt1_driver.sv
`include agnt1_mon.sv
`include agnt1_seqr.sv
`include agnt1_agent.sv
endpackage
