package agnt_pkg;
  import uvm_pkg::*;
  import struct_pkg::*;
  `include "uvm_macros.svh"
  `include "axi_narrow_seq_item.sv"
  `include "axi_narrow_driver.sv"
  `include "axi_narrow_mon.sv"
  `include "axi_narrow_seqr.sv"
  `include "axi_narrow_agent.sv"
  `include "axi_narrow_sequence.sv"
  `include "axi_wide_seq_item.sv"
  `include "axi_wide_driver.sv"
  `include "axi_wide_mon.sv"
  `include "axi_wide_seqr.sv"
  `include "axi_wide_agent.sv"
  `include "axi_wide_sequence.sv"
endpackage
