package agnt2_pkg;
`include agnt2_seq_item.sv
`include agnt2_driver.sv
`include agnt2_mon.sv
`include agnt2_seqr.sv
`include agnt2_agent.sv
endpackage
