package struct_pkg;
  `include "axi_narrow_struct.sv"
  `include "axi_wide_struct.sv"
endpackage
