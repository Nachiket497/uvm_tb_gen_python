interface dut_intf;
endinterface
