package sequence_pkg;
`include  "axi_narrow_sequence.sv"
 `include  "axi_wide_sequence.sv"
 endpackage
