interface intf_name;


endinterface
