module dut_top_wrapper(
    clk_reset_if        clk_reset_intf
       ,axi_narrow_intf axi_narrow_intf_h
       ,axi_wide_intf axi_wide_intf_h
   );

endmodule
