package dut_agnt_pkg;
`include "agnt1_pkg.sv"
import agnt1_pkg::*;
`include "agnt2_pkg.sv"
import agnt2_pkg::*;
endpackage
