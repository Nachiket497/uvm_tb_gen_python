package axi_wide_pkg;
  `include "axi_wide_seq_item.sv"
  `include "axi_wide_driver.sv"
  `include "axi_wide_mon.sv"
  `include "axi_wide_seqr.sv"
  `include "axi_wide_agent.sv"
  `include "axi_wide_sequence.sv"
endpackage
