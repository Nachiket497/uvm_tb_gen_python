package axi_narrow_pkg;
  `include "axi_narrow_seq_item.sv"
  `include "axi_narrow_driver.sv"
  `include "axi_narrow_mon.sv"
  `include "axi_narrow_seqr.sv"
  `include "axi_narrow_agent.sv"
  `include "axi_narrow_sequence.sv"
endpackage
